module parking_system (
    
);
    
endmodule